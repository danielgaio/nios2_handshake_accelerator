-- Qsys_handshake_tb.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Qsys_handshake_tb is
end entity Qsys_handshake_tb;

architecture rtl of Qsys_handshake_tb is
	component Qsys_handshake is
		port (
			clk_clk       : in std_logic := 'X'; -- clk
			reset_reset_n : in std_logic := 'X'  -- reset_n
		);
	end component Qsys_handshake;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal qsys_handshake_inst_clk_bfm_clk_clk       : std_logic; -- Qsys_handshake_inst_clk_bfm:clk -> [Qsys_handshake_inst:clk_clk, Qsys_handshake_inst_reset_bfm:clk]
	signal qsys_handshake_inst_reset_bfm_reset_reset : std_logic; -- Qsys_handshake_inst_reset_bfm:reset -> Qsys_handshake_inst:reset_reset_n

begin

	qsys_handshake_inst : component Qsys_handshake
		port map (
			clk_clk       => qsys_handshake_inst_clk_bfm_clk_clk,       --   clk.clk
			reset_reset_n => qsys_handshake_inst_reset_bfm_reset_reset  -- reset.reset_n
		);

	qsys_handshake_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => qsys_handshake_inst_clk_bfm_clk_clk  -- clk.clk
		);

	qsys_handshake_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => qsys_handshake_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => qsys_handshake_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of Qsys_handshake_tb
